library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity Registrador is
generic(
	   DATA_WIDTH : natural := 64);
port ( i_RESET : in  std_logic;  -- clear/reset
       i_CLK   : in  std_logic;  -- clock
       i_ENA   : in  std_logic;  -- enable    
       i_D     : in  std_logic_vector(DATA_WIDTH-1 downto 0);  -- data input
       o_Q     : out std_logic_vector(DATA_WIDTH-1 downto 0)); -- data output
end Registrador;


architecture arch_Reg of Registrador is
	signal w_EX_SIGNAL : std_logic_vector(DATA_WIDTH-1 downto 0);
begin
  process(i_RESET,i_CLK) 
  begin
    if (i_RESET ='1') then
      o_Q <= (others =>'0');
	elsif (rising_edge(i_CLK)) then
      if (i_ENA = '1') then
         o_Q <= i_D;
      end if;
    end if;
  end process;
end arch_Reg;